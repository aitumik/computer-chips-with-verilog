module main;

  initial
    begin
      $display("Learning Verilog is easy with me");
      $finish;
    end
endmodule
