module data_selector(
  input A,
  input B,
  input SEL,
  output Q
);

endmodule
